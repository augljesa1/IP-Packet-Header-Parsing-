LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY IPv4_PARSING_HEADER_testbench IS
END IPv4_PARSING_HEADER_testbench;

ARCHITECTURE arch_IPv4_PARSING_HEADER_testbench OF IPv4_PARSING_HEADER_testbench IS
COMPONENT IPv4_PARSING_HEADER IS
	PORT (
		PACKET : IN  STD_LOGIC_VECTOR(511 DOWNTO 0);
		MAC_SRC: OUT  STD_LOGIC_VECTOR(47 DOWNTO 0);
	   MAC_DST: OUT  STD_LOGIC_VECTOR(47 DOWNTO 0);
		MAC_BROADCAST : OUT  STD_LOGIC;
	   IPv4_VALID : OUT STD_LOGIC;
	   IPv4_SRC : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	   IPv4_DST : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	   IPv4_CLASS_A : OUT STD_LOGIC;
	   IPv4_CLASS_B : OUT STD_LOGIC;
	   IPv4_CLASS_C : OUT STD_LOGIC;
	   IPv4_BROADCAST : OUT STD_LOGIC;
	   IPv4_TTL: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

SIGNAL s_PACKET : STD_LOGIC_VECTOR(511 DOWNTO 0);
SIGNAL s_MAC_SRC, s_MAC_DST : STD_LOGIC_VECTOR(47 DOWNTO 0);
SIGNAL s_IPv4_SRC, s_IPv4_DST : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL s_IPv4_TTL : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL s_MAC_BROADCAST, s_IPv4_VALID, s_IPv4_CLASS_A, s_IPv4_CLASS_B, s_IPv4_CLASS_C, s_IPv4_BROADCAST : STD_LOGIC;

BEGIN
uut: IPv4_PARSING_HEADER
PORT MAP (
	PACKET => s_PACKET,
	MAC_SRC => s_MAC_SRC,
	MAC_DST => s_MAC_DST,
	MAC_BROADCAST => s_MAC_BROADCAST,
	IPv4_VALID => s_IPv4_VALID,
	IPv4_SRC => s_IPv4_SRC,
	IPv4_DST => s_IPv4_DST,
	IPv4_CLASS_A => s_IPv4_CLASS_A,
	IPv4_CLASS_B => s_IPv4_CLASS_B,
	IPv4_CLASS_C => s_IPv4_CLASS_C,
	IPv4_BROADCAST => s_IPv4_BROADCAST,
	IPv4_TTL => s_IPv4_TTL
	);
	
stim: PROCESS
BEGIN
  
  s_PACKET <= "11000110101001011001000110010100110101010100010111110100101101011001000110010100110101010100010010101010101100101000110101001011001000110001010011010101010001010101011101010101110001101010010100110000110010011101010101000100010101100101000111111111111111111111111111111111110101010110010101010111010101011100011010100101000100011001010011010101010111010101011101010101110001101010010100010001100101001101010101001101010101110101010111000110101001010001000110010100110101010100010101010111010101011100011010100101";

  WAIT;
END PROCESS;
verif: PROCESS

BEGIN
  --provjera izlaza za paket(checksum, IP i MAC adrese, IP broadcast, TTL)
  --WAIT FOR 10 ns;
  ASSERT (s_MAC_DST = "110001101010010110010001100101001101010101000101") REPORT "Greska 1" SEVERITY error;
  ASSERT (s_MAC_SRC = "111101001011010110010001100101001101010101000100") REPORT "Greska 2" SEVERITY error;
  ASSERT (s_IPV4_SRC = "11010101010001000101011001010001") REPORT "Greska 3" SEVERITY error;
  ASSERT (s_IPV4_DST = "11111111111111111111111111111111") REPORT "Greska 4" SEVERITY error;
  ASSERT (s_MAC_BROADCAST = '1') REPORT "Greska 5" SEVERITY error;
  ASSERT (s_IPv4_BROADCAST = '1') REPORT "Greska 6" SEVERITY error; 
  ASSERT (s_IPv4_CLASS_A = '1') REPORT "Greska 7" SEVERITY error;
  ASSERT (s_IPv4_CLASS_B = '1') REPORT "Greska 8" SEVERITY error; 
  ASSERT (s_IPv4_CLASS_C = '1') REPORT "Greska 9" SEVERITY error; 
  ASSERT (s_IPv4_TTL = "11000110") REPORT "Greska 10" SEVERITY error;
  ASSERT (s_IPv4_VALID = '1') REPORT "Greska 11" SEVERITY error;
   
  WAIT;

 END PROCESS;
END ARCHITECTURE;