LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY IPv4_PARSING_HEADER3_testbench IS
END IPv4_PARSING_HEADER3_testbench;

ARCHITECTURE arch_IPv4_PARSING_HEADER3_testbench OF IPv4_PARSING_HEADER3_testbench IS
COMPONENT IPv4_PARSING_HEADER IS
	PORT (
		PACKET : IN  STD_LOGIC_VECTOR(511 DOWNTO 0);
		MAC_SRC: OUT  STD_LOGIC_VECTOR(47 DOWNTO 0);
	   MAC_DST: OUT  STD_LOGIC_VECTOR(47 DOWNTO 0);
		MAC_BROADCAST : OUT  STD_LOGIC;
	   IPv4_VALID : OUT STD_LOGIC;
	   IPv4_SRC : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	   IPv4_DST : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	   IPv4_CLASS_A : OUT STD_LOGIC;
	   IPv4_CLASS_B : OUT STD_LOGIC;
	   IPv4_CLASS_C : OUT STD_LOGIC;
	   IPv4_BROADCAST : OUT STD_LOGIC;
	   IPv4_TTL: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

SIGNAL s_PACKET : STD_LOGIC_VECTOR(511 DOWNTO 0);
SIGNAL s_MAC_SRC, s_MAC_DST : STD_LOGIC_VECTOR(47 DOWNTO 0);
SIGNAL s_IPv4_SRC, s_IPv4_DST : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL s_IPv4_TTL : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL s_MAC_BROADCAST, s_IPv4_VALID, s_IPv4_CLASS_A, s_IPv4_CLASS_B, s_IPv4_CLASS_C, s_IPv4_BROADCAST : STD_LOGIC;

BEGIN
uut: IPv4_PARSING_HEADER
PORT MAP (
	PACKET => s_PACKET,
	MAC_SRC => s_MAC_SRC,
	MAC_DST => s_MAC_DST,
	MAC_BROADCAST => s_MAC_BROADCAST,
	IPv4_VALID => s_IPv4_VALID,
	IPv4_SRC => s_IPv4_SRC,
	IPv4_DST => s_IPv4_DST,
	IPv4_CLASS_A => s_IPv4_CLASS_A,
	IPv4_CLASS_B => s_IPv4_CLASS_B,
	IPv4_CLASS_C => s_IPv4_CLASS_C,
	IPv4_BROADCAST => s_IPv4_BROADCAST,
	IPv4_TTL => s_IPv4_TTL
	);
stim: PROCESS
BEGIN
  
	s_PACKET <= "01010101101011101110101011101011010111011101011110101001010001011110101001010101000101010101111101010101011001011000110101001011011010100101010111000101001001101001101001101011101001010101010101010000001010010010011100101100101100010011010011001010101010101010101010101010101010101100101010101110101010111000110101001010001000110010100110101010101110101010111010101011100011010100101000100011001010011010101010011010101011101010101110001101011001010001000110010100110101010100010101010111010101011100011010100101";
          

  WAIT;
END PROCESS;
verif: PROCESS

BEGIN
  --provjera izlaza za prvi paket3(checksum, IP i MAC adrese, IP verzija C, TTL)
  WAIT FOR 10 ns;
  ASSERT (s_MAC_DST = "010101011010111011101010111010110101110111010111") REPORT "Greska 1" SEVERITY error; 
  ASSERT (s_MAC_SRC = "101010010100010111101010010101010001010101011111") REPORT "Greska 2" SEVERITY error;  
  ASSERT (s_IPV4_SRC = "00100111001011001011000100110100") REPORT "Greska 3" SEVERITY error; 
  ASSERT (s_IPV4_DST = "11001010101010101010101010101010") REPORT "Greska 4" SEVERITY error;  
  ASSERT (s_MAC_BROADCAST = '1') REPORT "Greska 5" SEVERITY error; 
  ASSERT (s_IPv4_BROADCAST = '1') REPORT "Greska 6" SEVERITY error; 
  ASSERT (s_IPv4_CLASS_A = '1') REPORT "Greska 7" SEVERITY error;
  ASSERT (s_IPv4_CLASS_B = '1') REPORT "Greska 8" SEVERITY error;
  ASSERT (s_IPv4_CLASS_C = '1') REPORT "Greska 9" SEVERITY error; 
  ASSERT (s_IPv4_TTL = "10100101") REPORT "Greska 10" SEVERITY error; 
  ASSERT (s_IPv4_VALID = '1') REPORT "Greska 11" SEVERITY error;  
  
  WAIT;

 END PROCESS;
END ARCHITECTURE;
	


